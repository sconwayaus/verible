module tabs;
	int a; // tabs bad!
endmodule
