// Expects module port 'hello_world' to be lower_snakecase with _i suffix
module port_name_style(input bit hello_world);  // verilog_lint: waive port-name-suffix
endmodule
