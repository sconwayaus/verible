// Expects module port 'hello_world' to follow end with _i
module port_name_suffix(input bit hello_world);  // verilog_lint: waive port-name-style
endmodule
