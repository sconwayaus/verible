// Expects signal 'helloWorld' to follow lower_snake_case naming convention.
module signal_name_style();
    logic helloWorld;
endmodule
